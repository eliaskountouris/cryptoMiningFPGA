module sha256
(
    input logic [31:letters
);

endmodule
