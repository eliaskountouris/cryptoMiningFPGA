../../desigin/sha256/sha256.sv